library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Font_ROM is
	port(
		addr: in std_logic_vector(8 downto 0);
		data: out std_logic_vector(0 to 19)
	);
end Font_ROM;

architecture content of Font_ROM is
	type rom_type is array(0 to 191) of std_logic_vector(19 downto 0);
	
	constant FONT: rom_type :=
	(
		-- 0
		"00000001111111000000", --        #######      
		"00000101111111010000", --      # ####### #    
		"00000101111111011000", --      # ####### ##   
		"00001101111111011000", --     ## ####### ##   
		"00011100111111011100", --    ###  ###### ###  
		"00011100000000011110", --    ###         #### 
		"00111100000000011111", --   ####         #####
		"01111100000000011111", --  #####         #####
		"01111100000000011111", --  #####         #####
		"00000000000000000000", --                     
		"11111100000000011111", -- ######         #####
		"11111100000000011111", -- ######         #####
		"11111100000000011111", -- ######         #####
		"11111100000000011111", -- ######         #####
		"11111100000000011111", -- ######         #####
		"11111100000000011111", -- ######         #####
		"11111100000000011111", -- ######         #####
		"11111100000000011111", -- ######         #####
		"11111100000000011111", -- ######         #####
		"00000000000000000000", --                     
		"01111100111111011111", --  #####  ###### #####
		"01111101111111011111", --  ##### ####### #####
		"01111101111111011111", --  ##### ####### #####
		"00111101111111011110", --   #### ####### #### 
		"00011101111111011110", --    ### ####### #### 
		"00011101111111011100", --    ### ####### ###  
		"00001101111111011000", --     ## ####### ##   
		"00000101111111010000", --      # ####### #    
		"00000001111111010000", --        ####### #    
		"00000001111111000000", --        #######      
		"00000000000000000000", --                     
		"00000000000000000000", --                     

		-- 1
		"00000001111111000000", --        #######      
		"00000101111111000000", --      # #######      
		"00000101111111000000", --      # #######      
		"00001101111111000000", --     ## #######      
		"00011101111111000000", --    ### #######      
		"00111101111111000000", --   #### #######      
		"00111101111111000000", --   #### #######      
		"01111101111111000000", --  ##### #######      
		"11111101111111000000", -- ###### #######      
		"11111100000000000000", -- ######              
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000000000000000000", --                     
		"00000001111110000000", --        ######       
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000001111111000000", --        #######      
		"00000000000000000000", --                     
		"00000000000000000000", --                     

		-- 2
		"11111011111100000000", -- ##### ######        
		"11111011111101100000", -- ##### ###### ##     
		"11111011111101100000", -- ##### ###### ##     
		"11111011111101110000", -- ##### ###### ###    
		"11111011111101111000", -- ##### ###### ####   
		"00000000000001111000", --              ####   
		"00000000000001111100", --              #####  
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000000000000", --                     
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111000000000000000", -- #####               
		"11111000000000000000", -- #####               
		"11111000000000000000", -- #####               
		"11111000000000000000", -- #####               
		"00000000000000000000", --                     
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"00000000000000000000", --                     
		"00000000000000000000", --                     

		-- 3
		"11111011111100000000", -- ##### ######        
		"11111011111101000000", -- ##### ###### #      
		"11111011111101100000", -- ##### ###### ##     
		"11111011111101100000", -- ##### ###### ##     
		"11110011111101110000", -- ####  ###### ###    
		"00000000000001111000", --              ####   
		"00000000000001111100", --              #####  
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000000000000", --                     
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11110011111101111111", -- ####  ###### #######
		"00000000000001111111", --              #######
		"00000000000001111111", --              #######
		"00000000000001111111", --              #######
		"00000000000001111111", --              #######
		"00000000000000000000", --                     
		"11111011111101111110", -- ##### ###### ###### 
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"00000000000000000000", --                     
		"00000000000000000000", --                     

		-- 4
		"11110000000000000000", -- ####                
		"11110000000001000000", -- ####         #      
		"11110000000001000000", -- ####         #      
		"11110000000001100000", -- ####         ##     
		"11110000000001110000", -- ####         ###    
		"11110000000001110000", -- ####         ###    
		"11110000000001111000", -- ####         ####   
		"11110000000001111100", -- ####         #####  
		"11110000000001111100", -- ####         #####  
		"00000000000000000000", --                     
		"11110011111101111110", -- ####  ###### ###### 
		"11110011111101111110", -- ####  ###### ###### 
		"11110011111101111110", -- ####  ###### ###### 
		"11110011111101111110", -- ####  ###### ###### 
		"11110011111101111110", -- ####  ###### ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000000000000", --                     
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000000000000", --                     
		"00000000000000000000", --                     

		-- 5
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111000000000000000", -- #####               
		"11111000000000000000", -- #####               
		"11111000000000000000", -- #####               
		"11111000000000000000", -- #####               
		"11111000000000000000", -- #####               
		"00000000000000000000", --                     
		"11111011111100000000", -- ##### ######        
		"11111011111101000000", -- ##### ###### #      
		"11111011111101100000", -- ##### ###### ##     
		"11111011111101110000", -- ##### ###### ###    
		"11111011111101111000", -- ##### ###### ####   
		"00000000000001111000", --              ####   
		"00000000000001111100", --              #####  
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000001111110", --              ###### 
		"00000000000000000000", --                     
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"11111011111101111111", -- ##### ###### #######
		"00000000000000000000", --                     
		"00000000000000000000"  --                     
	);
begin
	data <= FONT(conv_integer(addr));
end content;