package dlx_package is

	constant c_DLX_PC_WIDTH : integer := 10;
	constant c_DLX_WORD_WIDTH : integer := 32;

end package dlx_package;

package body dlx_package is

end package body dlx_package;